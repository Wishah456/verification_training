package pkg;
  //  Group: Typedefs
  typedef class animal;
  typedef class bird;

  //  Group: Parameters
  `include "animal.svh"
  `include "bird.svh"

endpackage
